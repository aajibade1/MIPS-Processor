`include "types_pkg.vh"

module test_fpga (
  input logic [3:0] KEY,
  output logic [6:0]HEX0
);
  import types_pkg::*;
  my_t myvalue;

  test DUT(
    .CLK (~KEY[3]),
    .nRST (KEY[0]),
    .down (~KEY[2]),
    .value (myvalue)
  );

  always_comb
  begin
    unique casez (myvalue)
      'h0: HEX0 = 7'b1000000;
      'h1: HEX0 = 7'b1111001;
      'h2: HEX0 = 7'b0100100;
      'h3: HEX0 = 7'b0110000;
      'h4: HEX0 = 7'b0011001;
      'h5: HEX0 = 7'b0010010;
      'h6: HEX0 = 7'b0000010;
      'h7: HEX0 = 7'b1111000;
      'h8: HEX0 = 7'b0000000;
      'h9: HEX0 = 7'b0010000;
      'ha: HEX0 = 7'b0001000;
      'hb: HEX0 = 7'b0000011;
      'hc: HEX0 = 7'b0100111;
      'hd: HEX0 = 7'b0100001;
      'he: HEX0 = 7'b0000110;
      'hf: HEX0 = 7'b0001110;
    endcase
  end
endmodule
