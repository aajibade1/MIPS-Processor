/*
  sample package
*/
`ifndef TYPES_PKG_VH
`define TYPES_PKG_VH
package types_pkg;
  typedef logic [3:0] my_t;
endpackage
`endif //TYPES_PKG_VH
